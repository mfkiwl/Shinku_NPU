module instr_ram #(parameter WIDTH = 32)
(
	input [31:0] d,
	input [31:0] addr,
	input clk, menable,
	output reg [31:0] q
);

	// Declare the RAM variable
	reg [31:0] ram[1024:0];
	
	initial begin
//	 integer i;
//    for(i=0;i<63;i=i+1)
//       ram[i]=0;
		ram[32'h00000000] = 32'h0000_0013; //  NOP(to wait to finish register load)
		ram[32'h00000004] = 32'h0000_6183; //	load 512bit,$512_3,0x0000_0000
		ram[32'h00000008] = 32'h0010_6203; //  load 512bit,$512_4,0x0000_0081
		ram[32'h0000000c] = 32'h0020_6283; //	load 512bit,$512_5,0x0000_0102	
		ram[32'h00000010] = 32'h0030_6303; //  load 512bit,$512_6,0x0000_0183
		ram[32'h00000014] = 32'h0040_6383; //  load 512bit,$512_7,0x0000_0204
		ram[32'h00000018] = 32'h0000_0013; //  NOP(to wait to finish register load)
		ram[32'h0000001c] = 32'h0000_0013; //  NOP(to wait to finish register load)
		ram[32'h00000020] = 32'h0000_0013; //  NOP(to wait to finish register load)
		ram[32'h00000024] = 32'h0000_00AB; //  NWL Load Network, $512_1
		ram[32'h00000028] = 32'h0030_F10B; //	NWAND $512_1,$512_3,$512_2
		ram[32'h0000002c] = 32'h0040_F08B; //  NWAND $512_1,$512_4,$512_1
		ram[32'h00000030] = 32'h0060_908B; //  NWSLL $512_1,$512_6,$512_1
		ram[32'h00000034] = 32'h0020_E08B; //  NWOR  $512_1,$512_2,$512_1
		ram[32'h00000038] = 32'h0050_E08B; //	NWOR  $512_1,$512_5,$512_1
      ram[32'h0000003c] = 32'h0070_808B; //	NWADD  $512_1,$512_7,$512_1
		ram[32'h00000040] = 32'h0010_102B; //	NWS Store Network, $512_1
		ram[32'h00000044] = 32'hFDDF_F06F; //	jmp PC-0x14

	end
		
	always @(negedge clk)
	begin
	// Write
		if (menable == 1) ram[addr] <= d;
	//read
		q <= ram[addr];		
	end
	

endmodule

module data_ram #(parameter WIDTH = 32)
(
	input [31:0] d,
//	input [511:0] d_512,
	input [31:0] addr,
//	input [2:0] rmode,wmode,
	input clk, menable,
	output reg [31:0] q
//	output reg [511:0] q_512
);

	// Declare the RAM variable
	reg [31:0] ram[4096:0];
	
		always @(negedge clk)
	begin
	// Write
		if (menable == 1) ram[addr] <= d;
	//read
		q <= ram[addr];		
	end

		 initial begin

        end

endmodule

module data_ram_1024 #(parameter WIDTH = 32)
(
	input [1047:0] d,
	input [31:0] addr,
	input clk, menable,
	output reg [1047:0] q
);

	// Declare the RAM variable
	reg [1047:0]ram[1024:0];
	
	initial begin
		//bitmask For HEADER(MAC address)
		ram[32'h0000_0000] <= 1048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF_FFFF_FF;
		
		//Bitmask for DATA 
		ram[32'h0000_0001] <= 1048'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000_0000_00;
		
		//VLAN header data
		ram[32'h0000_0002] <= 1048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002000018000000000000000000000000_0000_00;
		
		//DATA shift amount
		ram[32'h0000_0003] <= 1048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000020;

        //ADD DATA (1)
        ram[32'h0000_0004] <= 1048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000004;
	end
				
	always @(negedge clk)
	begin
	// Write
		if (menable == 1) ram[addr] <= d;
	//read
		q <= ram[addr];		
	end

endmodule

